/*
 * Shifter_tb.sv
 * Shawn Zhu
 * ECE552
 */
module Shifter_tb();
reg signed [15:0] Shift_In; 	// This is the input data to perform shift operation on
reg [3:0] Shift_Val; 	// Shift amount (used to shift the input data)
reg  [1:0] Mode; 	// To indicate 0=SLL or 1=SRA 
wire [15:0] Shift_Out; 	// Shifted output data

Shifter DUT(.Shift_Out(Shift_Out), .Shift_In(Shift_In), .Shift_Val(Shift_Val), .Mode(Mode));

logic [15:0] shift_check = 0;
logic [15:0] shift_res = 0;
logic [15:0] shift_out = 0;
initial begin
	$randomize;
	repeat(50) begin
		//set inputs to be random
		Shift_In = $random;
		Shift_Val = $random;
		Mode = $urandom_range(0, 2);
		
		// display inputs
		$display("Test Case %0d:", $time);
		$display("Input: %b, Shift Amount: %b, Mode: %b", Shift_In, Shift_Val, Mode);
		
		//generate the shift results
		if(Mode[1] && ~Mode[0]) begin
			shift_res = Shift_In >> Shift_Val;
			shift_out = Shift_In << 16 - Shift_Val;
			shift_check = shift_res | shift_out;
		end
		else if (Mode[1] && Mode[0]) begin
			$error("Unused Opcode");
		end
		else begin
			if(Mode[0]) shift_check = Shift_In >>> Shift_Val;
			else shift_check = Shift_In << Shift_Val;
		end
		
		#1
		$display("Result: %b", Shift_Out);
		
		//check if the shifter worked
		if(shift_check != Shift_Out) $error("TEST FAILED");
		else $display("TEST PASSED");
	end
end

endmodule
