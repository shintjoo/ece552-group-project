/*
 * PADDSB_tb.sv
 * Shawn Zhu
 * ECE552
 */
module PADDSB_tb ();
reg [15:0] A, B;
wire [15:0] Sum;

endmodule